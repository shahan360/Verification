// Code your testbench here
// or browse Examples
`include "uvm_macros.svh"
import uvm_pkg::*;

module top;
  initial begin
    `uvm_info("TESTTOP","My first UVM testbench!", UVM_NONE);
  end
  
endmodule  